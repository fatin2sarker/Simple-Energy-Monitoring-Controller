LIBRARY ieee;
USE ieee.std_logic_1164.all;
LIBRARY work;
ENTITY VHDL_polarity_control IS
       PORT  (
		       POLARITY_CNTRL,XOR_IN1,XOR_IN2,XOR_IN3,XOR_IN4 : IN STD_LOGIC; XOR_OUT1, XOR_OUT2, XOR_OUT3, XOR_OUT4 : OUT STD_LOGIC
				 );
END VHDL_polarity_control;

ARCHITECTURE simple_gates OF VHDL_polarity_control IS
BEGIN

XOR_OUT1 <= POLARITY_CNTRL XOR XOR_IN1;
XOR_OUT2 <= POLARITY_CNTRL XOR XOR_IN2;
XOR_OUT3 <= POLARITY_CNTRL XOR XOR_IN3;
XOR_OUT4 <= POLARITY_CNTRL XOR XOR_IN4;


END ARCHITECTURE simple_gates;